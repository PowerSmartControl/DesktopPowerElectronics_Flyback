** Profile: "Control-Temp"  [ C:\Documents and Settings\EGA\Escritorio\convertidor ac-dc-pspicefiles\control\temp.sim ] 

** Creating circuit file "Temp.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "E:/Hardware/OrCAD/Capture/PSpice/burr_brn.lib" 
* From [PSPICE NETLIST] section of E:\zOrCAD\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 80ms 0 .2ms 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Control.net" 


.END
